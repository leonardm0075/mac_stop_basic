`timescale 1ns / 1ps

module test_mac_stop_accum;
    //Test Case 1: Matrix A is 2x2 and matrix B is 2x2 --> M = 2, K = 2, N = 2 --> all prduct and accumulation values fall in the decimal range of 0-50
    //Test Case 2: Matrix A is 10x8 and matrix B is 8x5 --> M = 10, K = 8, N = 5 --> all prduct and accumulation values fall in the decimal range of 50-100
    //Test Case 3: Matrix A is 3x5 and matrix B is 5x5 --> M = 3, K = 5, N = 5 --> all prduct and accumulation values fall in the decimal range of 100-150

    // Parameters
    parameter M = 3;
    parameter K = 5;
    parameter N = 5;
    parameter DATA_WIDTH_INIT_MATRIX = 32;
    parameter DATA_WIDTH_RESULT_MATRIX = (DATA_WIDTH_INIT_MATRIX * 2 + $clog2(K));

    // Inputs
    logic clk;
    logic resetn;
    logic [(DATA_WIDTH_INIT_MATRIX*2)-1:0] product_reg;
    logic [$clog2(K)-1:0] matrix_a_col_addr_counter_reg, matrix_b_row_addr_counter_reg;
    logic [$clog2(M)-1:0] matrix_a_row_addr_counter_reg;
    logic [$clog2(N)-1:0] matrix_b_col_addr_counter_reg;
    logic mult_done_reg;

    // Outputs
    logic [DATA_WIDTH_RESULT_MATRIX-1:0] data_out_c;
    logic matrix_c_we;
    logic mac_done;
    logic [$clog2(M)-1:0] row_addr_c;
    logic [$clog2(N)-1:0] col_addr_c;

    // Instantiate the Unit Under Test (UUT)
    mac_stop #(
        .M(M),
        .K(K),
        .N(N),
        .DATA_WIDTH_INIT_MATRIX(DATA_WIDTH_INIT_MATRIX),
        .DATA_WIDTH_RESULT_MATRIX(DATA_WIDTH_RESULT_MATRIX)
    ) uut (
        .clk(clk),
        .resetn(resetn),
        .data_out_c(data_out_c),
        .matrix_c_we(matrix_c_we),
        .product_reg(product_reg),
        .matrix_a_col_addr_counter_reg(matrix_a_col_addr_counter_reg),
        .matrix_b_row_addr_counter_reg(matrix_b_row_addr_counter_reg),
        .matrix_a_row_addr_counter_reg(matrix_a_row_addr_counter_reg),
        .matrix_b_col_addr_counter_reg(matrix_b_col_addr_counter_reg),
        .mult_done_reg(mult_done_reg),
        .mac_done(mac_done),
        .row_addr_c(row_addr_c),
        .col_addr_c(col_addr_c)
    );

    logic [(M*N*K)-1:0][(DATA_WIDTH_INIT_MATRIX*2)-1:0] product_reg_array;
    logic [(M*N*K)-1:0][$clog2(K)-1:0] matrix_a_col_addr_counter_reg_array, matrix_b_row_addr_counter_reg_array;
    logic [(M*N*K)-1:0][$clog2(M)-1:0] matrix_a_row_addr_counter_reg_array;
    logic [(M*N*K)-1:0][$clog2(N)-1:0] matrix_b_col_addr_counter_reg_array;
    

    // Clock generation
    always #5 clk = ~clk;

    initial begin
        // Initialize Inputs
        clk = 0;
        resetn = 0;
        product_reg = 0;
        matrix_a_col_addr_counter_reg = 0;
        matrix_b_row_addr_counter_reg = 0;
        matrix_a_row_addr_counter_reg = 0;
        matrix_b_col_addr_counter_reg = 0;
        mult_done_reg = 0;

        //Test Case 1 values
        //product_reg_array = '{32, 18, 28, 15, 16, 6, 14, 5};
        //matrix_a_col_addr_counter_reg_array = '{1,0,1,0,1,0,1,0};
        //matrix_b_row_addr_counter_reg_array = '{1,0,1,0,1,0,1,0};
        //matrix_a_row_addr_counter_reg_array = '{1,1,1,1,0,0,0,0};
        //matrix_b_col_addr_counter_reg_array = '{1,1,0,0,1,1,0,0};

        //Test Case 2 values
        //product_reg_array = '{12, 4, 1, 16, 12, 9, 4, 2, 12, 3, 4, 16, 6, 6, 6, 2, 6, 3, 4, 16, 12, 6, 2, 2, 6, 1, 2, 16, 12, 12, 4, 1, 3, 1, 2, 12, 12, 12, 6, 4, 12, 4, 2, 12, 12, 6, 8, 2, 12, 3, 8, 12, 6, 4, 12, 2, 6, 3, 8, 12, 12, 4, 4, 2, 6, 1, 4, 12, 12, 8, 8, 1, 3, 1, 4, 9, 12, 8, 12, 4, 16, 4, 3, 8, 4, 12, 6, 8, 16, 3, 12, 8, 2, 8, 9, 8, 8, 3, 12, 8, 4, 8, 3, 8, 8, 1, 6, 8, 4, 16, 6, 4, 4, 1, 6, 6, 4, 16, 9, 16, 16, 12, 4, 12, 12, 9, 2, 2, 16, 9, 16, 12, 6, 6, 3, 2, 8, 9, 16, 12, 12, 6, 1, 2, 8, 3, 8, 12, 12, 12, 2, 1, 4, 3, 8, 9, 12, 12, 3, 4, 4, 8, 3, 16, 8, 12, 6, 4, 4, 6, 12, 16, 4, 8, 9, 4, 2, 6, 12, 16, 8, 8, 3, 4, 2, 2, 6, 16, 8, 16, 6, 2, 1, 2, 6, 12, 8, 16, 9, 8, 8, 16, 4, 16, 12, 6, 6, 8, 8, 12, 16, 16, 6, 4, 9, 8, 4, 12, 16, 16, 12, 4, 3, 8, 4, 4, 8, 16, 12, 8, 6, 4, 2, 4, 8, 12, 12, 8, 9, 16, 4, 8, 4, 8, 4, 12, 6, 8, 4, 6, 16, 8, 2, 8, 9, 8, 2, 6, 16, 8, 4, 8, 3, 8, 2, 2, 8, 8, 4, 16, 6, 4, 1, 2, 8, 6, 4, 16, 9, 16, 8, 12, 4, 12, 8, 12, 6, 6, 8, 9, 16, 12, 4, 8, 9, 6, 4, 9, 16, 12, 8, 8, 3, 6, 4, 3, 8, 12, 8, 16, 6, 3, 2, 3, 8, 9, 8, 16, 9, 12, 16, 12, 3, 16, 16, 6, 6, 2, 16, 9, 12, 16, 8, 4, 9, 2, 8, 9, 12, 16, 16, 4, 3, 2, 8, 3, 6, 16, 16, 8, 6, 1, 4, 3, 6, 12, 16, 8, 9, 4, 16, 16, 1, 16, 8, 9, 2, 8, 16, 12, 4, 16, 4, 6, 3, 8, 8, 12, 4, 16, 8, 6, 1, 8, 8, 4, 2, 16, 8, 12, 2, 4, 4, 4, 2, 12, 8, 12, 3, 16};
        //matrix_a_col_addr_counter_reg_array = '{7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0};
        //matrix_b_row_addr_counter_reg_array = '{7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0, 7, 6, 5, 4, 3, 2, 1, 0};
        //matrix_a_row_addr_counter_reg_array = '{9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 9, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 8, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 7, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 6, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 5, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0};
        //matrix_b_col_addr_counter_reg_array = '{4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0};

        //Test Case 3 Values
        product_reg_array = '{20, 18, 25, 24, 20, 24, 15, 25, 24, 20, 20, 18, 30, 20, 24, 20, 18, 25, 24, 20, 24, 15, 30, 20, 20, 15, 24, 20, 30, 20, 18, 20, 20, 30, 20, 15, 24, 24, 25, 24, 15, 24, 20, 30, 20, 18, 20, 24, 25, 20, 25, 24, 15, 24, 20, 30, 20, 15, 24, 20, 25, 24, 18, 20, 24, 25, 24, 15, 24, 20, 30, 20, 18, 20, 20};
        matrix_a_col_addr_counter_reg_array = '{4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0};
        matrix_b_row_addr_counter_reg_array = '{4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0, 4, 3, 2, 1, 0};
        matrix_a_row_addr_counter_reg_array = '{2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0, 0};
        matrix_b_col_addr_counter_reg_array = '{4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0, 4, 4, 4, 4, 4, 3, 3, 3, 3, 3, 2, 2, 2, 2, 2, 1, 1, 1, 1, 1, 0, 0, 0, 0, 0};



        // Reset the design
        #10; 
        resetn = 1;
        #10;

        for (int i=0; i<(M*N*K); i=i+1) begin
            mult_done_reg = 1;
            product_reg = product_reg_array[i];
            matrix_a_col_addr_counter_reg = matrix_a_col_addr_counter_reg_array[i];
            matrix_b_row_addr_counter_reg = matrix_b_row_addr_counter_reg_array[i];
            matrix_a_row_addr_counter_reg = matrix_a_row_addr_counter_reg_array[i];
            matrix_b_col_addr_counter_reg = matrix_b_col_addr_counter_reg_array[i];
            #5;
            if (matrix_c_we) begin
                $display("%0d: data_out_c = %d", i, data_out_c);
            end
            #5;

        end




        // Finish simulation
        #50 $finish;
    end

endmodule